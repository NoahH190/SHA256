module step_five (
    input [31:0]    i_w0, 
                    i_w1, 
                    i_w2, 
                    i_w3, 
                    i_w4, 
                    i_w5, 
                    i_w6, 
                    i_w7, 
                    i_w8, 
                    i_w9, 
                    i_w10, 
                    i_w11, 
                    i_w12, 
                    i_w13, 
                    i_w14, 
                    i_w15;

    input [31:0]    i_s00, 
                    i_s01, 
                    i_s02, 
                    i_s03, 
                    i_s04, 
                    i_s05, 
                    i_s06, 
                    i_s07, 
                    i_s08, 
                    i_s09, 
                    i_s010, 
                    i_s011, 
                    i_s012, 
                    i_s013, 
                    i_s014, 
                    i_s015;

    input [31:0]    i_s10, 
                    i_s11, 
                    i_s12, 
                    i_s13, 
                    i_s14, 
                    i_s15, 
                    i_s16, 
                    i_s17, 
                    i_s18, 
                    i_s19, 
                    i_s110, 
                    i_s111, 
                    i_s112, 
                    i_s113, 
                    i_s114, 
                    i_s115;

    output [31:0]   o_w16,
                    o_w17,
                    o_w18,
                    o_w19,
                    o_w20,
                    o_w21,
                    o_w22,
                    o_w23,
                    o_w24,
                    o_w25,
                    o_w26,
                    o_w27,
                    o_w28,
                    o_w29,
                    o_w30,
                    o_w31,
                    o_w32,
                    o_w33,
                    o_w34,
                    o_w35,
                    o_w36,
                    o_w37,
                    o_w38,
                    o_w39,
                    o_w40,
                    o_w41,
                    o_w42,
                    o_w43,
                    o_w44,
                    o_w45,
                    o_w46,
                    o_w47,
                    o_w48,
                    o_w49,
                    o_w50,
                    o_w51,
                    o_w52,
                    o_w53,
                    o_w54,
                    o_w55,
                    o_w56,
                    o_w57,
                    o_w58,
                    o_w59,
                    o_w60,
                    o_w61,
                    o_w62,
                    o_w63;
)

assign o_w16 = {i_w0,i_s00,i_w9,i_s10}