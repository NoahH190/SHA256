module step_two(
    input i_clk;
    input i_reset;
    input [31:0]    i_m0, 
                    i_m1, 
                    i_m2, 
                    i_m3, 
                    i_m4, 
                    i_m5, 
                    i_m6, 
                    i_m7, 
                    i_m8, 
                    i_m9, 
                    i_m10, 
                    i_m11, 
                    i_m12, 
                    i_m13, 
                    i_m14, 
                    i_m15;
    output [31:0]   o_w0, 
                    o_w1, 
                    o_w2, 
                    o_w3, 
                    o_w4, 
                    o_w5, 
                    o_w6, 
                    o_w7, 
                    o_w8, 
                    o_w9, 
                    o_w10, 
                    o_w11, 
                    o_w12, 
                    o_w13, 
                    o_w14, 
                    o_w15;
);



