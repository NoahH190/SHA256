module step_five (
    input [31:0]    i_w0, 
                    i_w1, 
                    i_w2, 
                    i_w3, 
                    i_w4, 
                    i_w5, 
                    i_w6, 
                    i_w7, 
                    i_w8, 
                    i_w9, 
                    i_w10, 
                    i_w11, 
                    i_w12, 
                    i_w13, 
                    i_w14, 
                    i_w15;

    output [31:0]   o_s00, 
                    o_s01, 
                    o_s02, 
                    o_s03, 
                    o_s04, 
                    o_s05, 
                    o_s06, 
                    o_s07, 
                    o_s08, 
                    o_s09, 
                    o_s010, 
                    o_s011, 
                    o_s012, 
                    o_s013, 
                    o_s014, 
                    o_s015;

    input [31:0]    o_s10, 
                    o_s11, 
                    o_s12, 
                    o_s13, 
                    o_s14, 
                    o_s15, 
                    o_s16, 
                    o_s17, 
                    o_s18, 
                    o_s19, 
                    o_s110, 
                    o_s111, 
                    o_s112, 
                    o_s113, 
                    o_s114, 
                    o_s115;

    output [31:0]   i_w16,
                    i_w17,
                    i_w18,
                    i_w19,
                    i_w20,
                    i_w21,
                    i_w22,
                    i_w23,
                    i_w24,
                    i_w25,
                    i_w26,
                    i_w27,
                    i_w28,
                    i_w29,
                    i_w30,
                    i_w31,
                    i_w32,
                    i_w33,
                    i_w34,
                    i_w35,
                    i_w36,
                    i_w37,
                    i_w38,
                    i_w39,
                    i_w40,
                    i_w41,
                    i_w42,
                    i_w43,
                    i_w44,
                    i_w45,
                    i_w46,
                    i_w47,
                    i_w48,
                    i_w49,
                    i_w50,
                    i_w51,
                    i_w52,
                    i_w53,
                    i_w54,
                    i_w55,
                    i_w56,
                    i_w57,
                    i_w58,
                    i_w59,
                    i_w60,
                    i_w61,
                    i_w62,
                    i_w63;
)

