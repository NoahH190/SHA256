module step_three(
    input i_clk;
    input i_reset;
    input [31:0]    i_w0, 
                    i_w1, 
                    i_w2, 
                    i_w3, 
                    i_w4, 
                    i_w5, 
                    i_w6, 
                    i_w7, 
                    i_w8, 
                    i_w9, 
                    i_w10, 
                    i_w11, 
                    i_w12, 
                    i_w13, 
                    i_w14, 
                    i_w15;
    output [31:0]   o_s00, 
                    o_s01, 
                    o_s02, 
                    o_s03, 
                    o_s04, 
                    o_s05, 
                    o_s06, 
                    o_s07, 
                    o_s08, 
                    o_s09, 
                    o_s010, 
                    o_s011, 
                    o_s012, 
                    o_s013, 
                    o_s014, 
                    o_s015;
);


