module step_three(
    input i_clk;
    input i_reset;
    input [31:0]    i_w0, 
                    i_w1, 
                    i_w2, 
                    i_w3, 
                    i_w4, 
                    i_w5, 
                    i_w6, 
                    i_w7, 
                    i_w8, 
                    i_w9, 
                    i_w10, 
                    i_w11, 
                    i_w12, 
                    i_w13, 
                    i_w14, 
                    i_w15;
    output [31:0]   o_s00, 
                    o_s01, 
                    o_s02, 
                    o_s03, 
                    o_s04, 
                    o_s05, 
                    o_s06, 
                    o_s07, 
                    o_s08, 
                    o_s09, 
                    o_s010, 
                    o_s011, 
                    o_s012, 
                    o_s013, 
                    o_s014, 
                    o_s015;
);

assign o_s00 = {i_w0[31:25], i_w0[24:0]}  ^ {i_w0[31:14], i_w0[13:0]}  ^ {3'b000, i_w0[28:0]};
assign o_s01 = {i_w1[31:25], i_w1[24:0]}  ^ {i_w1[31:14], i_w1[13:0]}  ^ {3'b000, i_w1[28:0]};
assign o_s02 = {i_w2[31:25], i_w2[24:0]}  ^ {i_w2[31:14], i_w2[13:0]}  ^ {3'b000, i_w2[28:0]};
assign o_s03 = {i_w3[31:25], i_w3[24:0]}  ^ {i_w3[31:14], i_w3[13:0]}  ^ {3'b000, i_w3[28:0]};
assign o_s04 = {i_w4[31:25], i_w4[24:0]}  ^ {i_w4[31:14], i_w4[13:0]}  ^ {3'b000, i_w4[28:0]};
assign o_s05 = {i_w5[31:25], i_w5[24:0]}  ^ {i_w5[31:14], i_w5[13:0]}  ^ {3'b000, i_w5[28:0]};
assign o_s06 = {i_w6[31:25], i_w6[24:0]}  ^ {i_w6[31:14], i_w6[13:0]}  ^ {3'b000, i_w6[28:0]};
assign o_s07 = {i_w7[31:25], i_w7[24:0]}  ^ {i_w7[31:14], i_w7[13:0]}  ^ {3'b000, i_w7[28:0]};
assign o_s08 = {i_w8[31:25], i_w8[24:0]}  ^ {i_w8[31:14], i_w8[13:0]}  ^ {3'b000, i_w8[28:0]};
assign o_s09 = {i_w9[31:25], i_w9[24:0]}  ^ {i_w9[31:14], i_w9[13:0]}  ^ {3'b000, i_w9[28:0]};
assign o_s010 = {i_w10[31:25], i_w10[24:0]} ^ {i_w10[31:14], i_w10[13:0]} ^ {3'b000, i_w10[28:0]};
assign o_s011 = {i_w11[31:25], i_w11[24:0]} ^ {i_w11[31:14], i_w11[13:0]} ^ {3'b000, i_w11[28:0]};
assign o_s012 = {i_w12[31:25], i_w12[24:0]} ^ {i_w12[31:14], i_w12[13:0]} ^ {3'b000, i_w12[28:0]};
assign o_s013 = {i_w13[31:25], i_w13[24:0]} ^ {i_w13[31:14], i_w13[13:0]} ^ {3'b000, i_w13[28:0]};
assign o_s014 = {i_w14[31:25], i_w14[24:0]} ^ {i_w14[31:14], i_w14[13:0]} ^ {3'b000, i_w14[28:0]};
assign o_s015 = {i_w15[31:25], i_w15[24:0]} ^ {i_w15[31:14], i_w15[13:0]} ^ {3'b000, i_w15[28:0]};

endmodule 